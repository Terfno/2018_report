** Profile: "SCHEMATIC1-exe3sim2"  [ W:\jkjs\exe3-schematic1-exe3sim2.sim ] 

** Creating circuit file "exe3-schematic1-exe3sim2.sim.cir" 
** WARNING: THIS AUTOMATICALLY GENERATED FILE MAY BE OVERWRITTEN BY SUBSEQUENT SIMULATIONS

*Libraries: 
* Local Libraries :
* From [PSPICE NETLIST] section of C:\Program Files\OrcadLite\PSpice\PSpice.ini file:
.lib "nom.lib" 

*Analysis directives: 
.TRAN  0 1.04 1.0 
.PROBE V(*) I(*) W(*) D(*) NOISE(*) 
.INC ".\exe3-SCHEMATIC1.net" 


.END
