** Profile: "SCHEMATIC1-exe3sim"  [ W:\jkjs\exe3-SCHEMATIC1-exe3sim.sim ] 

** Creating circuit file "exe3-SCHEMATIC1-exe3sim.sim.cir" 
** WARNING: THIS AUTOMATICALLY GENERATED FILE MAY BE OVERWRITTEN BY SUBSEQUENT SIMULATIONS

*Libraries: 
* Local Libraries :
* From [PSPICE NETLIST] section of C:\Program Files\OrcadLite\PSpice\PSpice.ini file:
.lib "nom.lib" 

*Analysis directives: 
.AC DEC 100 10 200
.PROBE V(*) I(*) W(*) D(*) NOISE(*) 
.INC ".\exe3-SCHEMATIC1.net" 


.END
